bind ptw ptw_prop
	#(
		.ASSERT_INPUTS (0)
	) u_ptw_sva(.*);