// The Clear BSD License
// Copyright (c) [2021] [The Trustees of Princeton University]
// All rights reserved.
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted for academic and research use only (subject to the 
// limitations in the disclaimer below) provided that the following conditions are met:
//     * Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
// 
//     * Redistributions in binary form must reproduce the above copyright
//     notice, this list of conditions and the following disclaimer in the
//     documentation and/or other materials provided with the distribution.
// 
//     * Neither the name of the copyright holder nor the names of its
//     contributors may be used to endorse or promote products derived from this
//     software without specific prior written permission.
// 
// NO EXPRESS OR IMPLIED LICENSES TO ANY PARTY'S PATENT RIGHTS ARE GRANTED BY
// THIS LICENSE. THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND
// CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
// PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
// CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,
// EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
// PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
// IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
// 
// This property file was autogenerated by AutoSVA on 2021-04-06
// to check the behavior of the original RTL module, whose interface is described below: 

/* verilator lint_off WIDTH */

module ptw_prop
 import ariane_pkg::*; #(
		parameter ASSERT_INPUTS = 0,
		parameter int ASID_WIDTH = 1,
		parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
		input  logic                    clk_i,                  // Clock
		input  logic                    rst_ni,                 // Asynchronous reset active low
		input  logic                    flush_i,                // flush everything, we need to do this because
		// actually everything we do is speculative at this stage
		// e.g.: there could be a CSR instruction that changes everything
		input  logic                    ptw_active_o, //output
		input  logic                    walking_instr_o,        // set when walking for TLB //output
		input  logic                    ptw_error_o,            // set when an error occurred //output
		input  logic                    ptw_access_exception_o, // set when an PMP access exception occured //output
		input  logic                    enable_translation_i,   // CSRs indicate to enable SV39
		input  logic                    en_ld_st_translation_i, // enable virtual memory translation for load/stores
		
		input  logic                    lsu_is_store_i,         // this translation was triggered by a store
		// PTW memory interface
		input  dcache_req_o_t           req_port_i,
		input  dcache_req_i_t           req_port_o, //output
		
		
		// to TLBs, update logic
		input  tlb_update_t             itlb_update_o, //output
		input  tlb_update_t             dtlb_update_o, //output
		
		input  logic [riscv::VLEN-1:0]  update_vaddr_o, //output
		
		input  logic [ASID_WIDTH-1:0]   asid_i,
		// from TLBs
		// did we miss?
		input  logic                    itlb_access_i,
		input  logic                    itlb_hit_i,
		input  logic [riscv::VLEN-1:0]  itlb_vaddr_i,
		
		input  logic                    dtlb_access_i,
		input  logic                    dtlb_hit_i,
		input  logic [riscv::VLEN-1:0]  dtlb_vaddr_i,
		// from CSR file
		input  logic [riscv::PPNW-1:0]  satp_ppn_i, // ppn from satp
		input  logic                    mxr_i,
		// Performance counters
		input  logic                    itlb_miss_o, //output
		input  logic                    dtlb_miss_o, //output
		// PMP
		
		input  riscv::pmpcfg_t [15:0]   pmpcfg_i,
		input  logic [15:0][53:0]       pmpaddr_i,
		input  logic [riscv::PLEN-1:0]  bad_paddr_o //output
		
	);

//==============================================================================
// Local Parameters
//==============================================================================

genvar j;
default clocking cb @(posedge clk_i);
endclocking
default disable iff (!rst_ni);

// Re-defined wires 
wire ptw_req_val;
wire ptw_req_rdy;
wire ptw_res_val;
wire itlb_iface_active;
wire itlb_val;
wire itlb_rdy;
wire [riscv::VLEN-1:0] itlb_stable;
wire [riscv::VLEN-1:0] itlb_data;
wire itlb_update_val;
wire [riscv::VLEN-1:0] itlb_update_data;
wire dtlb_iface_active;
wire dtlb_val;
wire dtlb_rdy;
wire [riscv::VLEN-1:0] dtlb_stable;
wire [riscv::VLEN-1:0] dtlb_data;
wire dtlb_update_val;
wire [riscv::VLEN-1:0] dtlb_update_data;

// Symbolics and Handshake signals
wire itlb_update_hsk = itlb_update_val;
wire itlb_hsk = itlb_val && itlb_rdy;
wire ptw_res_hsk = ptw_res_val;
wire ptw_req_hsk = ptw_req_val && ptw_req_rdy;
wire dtlb_update_hsk = dtlb_update_val;
wire dtlb_hsk = dtlb_val && dtlb_rdy;

//==============================================================================
// Modeling
//==============================================================================

// Modeling incoming request for itlb_iface
// Generate sampling signals and model
reg [3:0] itlb_iface_transid_sampled;
wire itlb_iface_transid_set = itlb_hsk;
wire itlb_iface_transid_response = itlb_update_hsk;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		itlb_iface_transid_sampled <= '0;
	end else if (itlb_iface_transid_set || itlb_iface_transid_response ) begin
		itlb_iface_transid_sampled <= itlb_iface_transid_sampled + itlb_iface_transid_set - itlb_iface_transid_response;
	end
end
co__itlb_iface_transid_sampled: cover property (|itlb_iface_transid_sampled);
if (ASSERT_INPUTS) begin
	as__itlb_iface_transid_sample_no_overflow: assert property (itlb_iface_transid_sampled != '1 || !itlb_iface_transid_set);
end else begin
	am__itlb_iface_transid_sample_no_overflow: assume property (itlb_iface_transid_sampled != '1 || !itlb_iface_transid_set);
end

as__itlb_iface_transid_active: assert property (itlb_iface_transid_sampled > 0 |-> itlb_iface_active);

// Assume payload is stable and valid is non-dropping
if (ASSERT_INPUTS) begin
	as__itlb_iface_transid_stability: assert property (itlb_val && !itlb_rdy |=> itlb_val && $stable(itlb_stable) );
end else begin
	am__itlb_iface_transid_stability: assume property (itlb_val && !itlb_rdy |=> itlb_val && $stable(itlb_stable) );
end

// Assert that if valid eventually ready or dropped valid
as__itlb_iface_transid_hsk_or_drop: assert property (itlb_val |-> s_eventually(!itlb_val || itlb_rdy));
// Assert that every request has a response and that every reponse has a request
as__itlb_iface_transid_eventual_response: assert property (itlb_iface_transid_set |-> s_eventually(itlb_update_val));
as__itlb_iface_transid_was_a_request: assert property (itlb_iface_transid_response |-> itlb_iface_transid_set || itlb_iface_transid_sampled);


// Modeling data integrity for itlb_iface_transid
reg [riscv::VLEN-1:0] itlb_iface_transid_data_model;
always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		itlb_iface_transid_data_model <= '0;
	end else if (itlb_iface_transid_set) begin
		itlb_iface_transid_data_model <= itlb_data;
	end
end

as__itlb_iface_transid_data_integrity: assert property (itlb_iface_transid_sampled && itlb_update_hsk |-> (itlb_update_data == itlb_iface_transid_data_model));

// Modeling outstanding request for ptw_req
reg [1-1:0] ptw_req_outstanding_req_r;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		ptw_req_outstanding_req_r <= '0;
	end else begin
		if (ptw_req_hsk) begin
			ptw_req_outstanding_req_r <= 1'b1;
		end
		if (ptw_res_hsk) begin
			ptw_req_outstanding_req_r <= 1'b0;
		end
	end
end


generate
if (ASSERT_INPUTS) begin : ptw_req_gen
	as__ptw_req1: assert property (!ptw_req_outstanding_req_r |-> !(ptw_res_hsk));
	as__ptw_req2: assert property (ptw_req_outstanding_req_r |-> s_eventually(ptw_res_hsk));
end else begin : ptw_req_else_gen
	am__ptw_req_fairness: assume property (ptw_req_val |-> s_eventually(ptw_req_rdy));
	for ( j = 0; j < 1; j = j + 1) begin : ptw_req_for_gen
		co__ptw_req: cover property (ptw_req_outstanding_req_r[j]);
		am__ptw_req1: assume property (!ptw_req_outstanding_req_r[j] |-> !(ptw_res_val));
		am__ptw_req2: assume property (ptw_req_outstanding_req_r[j] |-> s_eventually(ptw_res_val));
	end
end
endgenerate

// Modeling incoming request for dtlb_iface
// Generate sampling signals and model
reg [3:0] dtlb_iface_transid_sampled;
wire dtlb_iface_transid_set = dtlb_hsk;
wire dtlb_iface_transid_response = dtlb_update_hsk;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		dtlb_iface_transid_sampled <= '0;
	end else if (dtlb_iface_transid_set || dtlb_iface_transid_response ) begin
		dtlb_iface_transid_sampled <= dtlb_iface_transid_sampled + dtlb_iface_transid_set - dtlb_iface_transid_response;
	end
end
co__dtlb_iface_transid_sampled: cover property (|dtlb_iface_transid_sampled);
if (ASSERT_INPUTS) begin
	as__dtlb_iface_transid_sample_no_overflow: assert property (dtlb_iface_transid_sampled != '1 || !dtlb_iface_transid_set);
end else begin
	am__dtlb_iface_transid_sample_no_overflow: assume property (dtlb_iface_transid_sampled != '1 || !dtlb_iface_transid_set);
end

as__dtlb_iface_transid_active: assert property (dtlb_iface_transid_sampled > 0 |-> dtlb_iface_active);

// Assume payload is stable and valid is non-dropping
if (ASSERT_INPUTS) begin
	as__dtlb_iface_transid_stability: assert property (dtlb_val && !dtlb_rdy |=> dtlb_val && $stable(dtlb_stable) );
end else begin
	am__dtlb_iface_transid_stability: assume property (dtlb_val && !dtlb_rdy |=> dtlb_val && $stable(dtlb_stable) );
end

// Assert that if valid eventually ready or dropped valid
as__dtlb_iface_transid_hsk_or_drop: assert property (dtlb_val |-> s_eventually(!dtlb_val || dtlb_rdy));
// Assert that every request has a response and that every reponse has a request
as__dtlb_iface_transid_eventual_response: assert property (dtlb_iface_transid_set |-> s_eventually(dtlb_update_val));
as__dtlb_iface_transid_was_a_request: assert property (dtlb_iface_transid_response |-> dtlb_iface_transid_set || dtlb_iface_transid_sampled);


// Modeling data integrity for dtlb_iface_transid
reg [riscv::VLEN-1:0] dtlb_iface_transid_data_model;
always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		dtlb_iface_transid_data_model <= '0;
	end else if (dtlb_iface_transid_set) begin
		dtlb_iface_transid_data_model <= dtlb_data;
	end
end

as__dtlb_iface_transid_data_integrity: assert property (dtlb_iface_transid_sampled && dtlb_update_hsk |-> (dtlb_update_data == dtlb_iface_transid_data_model));

assign ptw_req_val = req_port_o.data_req;
assign dtlb_data = dtlb_vaddr_i;
assign itlb_update_val = itlb_update_o.valid || walking_instr_o && (ptw_access_exception_o || ptw_error_o || ptw_active_o && flush_i);
assign dtlb_update_val = dtlb_update_o.valid || !walking_instr_o && (ptw_access_exception_o || ptw_error_o || ptw_active_o && flush_i);
assign dtlb_val = en_ld_st_translation_i & dtlb_access_i & ~dtlb_hit_i & !flush_i;
assign dtlb_iface_active = ptw_active_o;
assign itlb_stable = itlb_vaddr_i;
assign dtlb_stable = dtlb_vaddr_i;
assign itlb_val = enable_translation_i & itlb_access_i & ~itlb_hit_i & ~dtlb_access_i & !flush_i;
assign ptw_req_rdy = req_port_i.data_gnt;
assign itlb_rdy = !ptw_active_o;
assign dtlb_rdy = !ptw_active_o;
assign dtlb_update_data = update_vaddr_o;
assign itlb_update_data = update_vaddr_o;
assign itlb_data = itlb_vaddr_i;
assign itlb_iface_active = ptw_active_o;
assign ptw_res_val = req_port_i.data_rvalid;

//X PROPAGATION ASSERTIONS
`ifdef XPROP
	 as__no_x_dtlb_update_val: assert property(!$isunknown(dtlb_update_val));
	 as__no_x_dtlb_update_data: assert property(dtlb_update_val |-> !$isunknown(dtlb_update_data));
	 as__no_x_dtlb_val: assert property(!$isunknown(dtlb_val));
	 as__no_x_dtlb_data: assert property(dtlb_val |-> !$isunknown(dtlb_data));
	 as__no_x_dtlb_stable: assert property(dtlb_val |-> !$isunknown(dtlb_stable));
	 as__no_x_itlb_update_val: assert property(!$isunknown(itlb_update_val));
	 as__no_x_itlb_update_data: assert property(itlb_update_val |-> !$isunknown(itlb_update_data));
	 as__no_x_itlb_val: assert property(!$isunknown(itlb_val));
	 as__no_x_itlb_stable: assert property(itlb_val |-> !$isunknown(itlb_stable));
	 as__no_x_itlb_data: assert property(itlb_val |-> !$isunknown(itlb_data));
`endif

//====DESIGNER-ADDED-SVA====//
am__1 : assume property (enable_translation_i);
am__2 : assume property (!flush_i);
endmodule