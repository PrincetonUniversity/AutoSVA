// The Clear BSD License
// Copyright (c) [2021] [The Trustees of Princeton University]
// All rights reserved.
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted for academic and research use only (subject to the 
// limitations in the disclaimer below) provided that the following conditions are met:
//     * Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
// 
//     * Redistributions in binary form must reproduce the above copyright
//     notice, this list of conditions and the following disclaimer in the
//     documentation and/or other materials provided with the distribution.
// 
//     * Neither the name of the copyright holder nor the names of its
//     contributors may be used to endorse or promote products derived from this
//     software without specific prior written permission.
// 
// NO EXPRESS OR IMPLIED LICENSES TO ANY PARTY'S PATENT RIGHTS ARE GRANTED BY
// THIS LICENSE. THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND
// CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
// PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
// CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,
// EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
// PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
// IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
// 
// This property file was autogenerated by AutoSVA on 2021-04-06
// to check the behavior of the original RTL module, whose interface is described below: 

// Author: Florian Zaruba, ETH Zurich
// Date: 19/04/2017
// Description: Memory Management Unit for Ariane, contains TLB and
//              address translation unit. SV39 as defined in RISC-V
//              privilege specification 1.11-WIP


module mmu_prop
 import ariane_pkg::*; #(
		parameter ASSERT_INPUTS = 0,
		parameter INSTR_TLB_ENTRIES     = 4,
		parameter DATA_TLB_ENTRIES      = 4,
		parameter ASID_WIDTH            = 1,
		parameter ariane_pkg::ariane_cfg_t ArianeCfg = 0//ariane_pkg::ArianeDefaultConfig
) (
		input  logic                            clk_i,
		input  logic                            rst_ni,
		input  logic                            flush_i,
		input  logic                            enable_translation_i,
		input  logic                            en_ld_st_translation_i,   // enable virtual memory translation for load/stores
		
		
		// IF interface
		input  icache_areq_o_t                  icache_areq_i,
		input  icache_areq_i_t                  icache_areq_o, //output
		
		// LSU interface
		// this is a more minimalistic interface because the actual addressing logic is handled
		// in the LSU as we distinguish load and stores, what we do here is simple address translation
		input  exception_t                      misaligned_ex_i,
		input  logic                            lsu_req_i,        // request address translation
		input  logic [riscv::VLEN-1:0]          lsu_vaddr_i,      // virtual address in
		input  logic                            lsu_is_store_i,   // the translation is requested by a store
		// if we need to walk the page table we can't grant in the same cycle
		// Cycle 0
		input  logic                            lsu_dtlb_hit_o,   // sent in the same cycle as the request if translation hits in the DTLB //output
		input  logic [riscv::PLEN-13:0]         lsu_dtlb_ppn_o,   // ppn (send same cycle as hit) //output
		// Cycle 1
		input  logic                            lsu_valid_o,      // translation is valid //output
		input  logic [riscv::PLEN-1:0]          lsu_paddr_o,      // translated address //output
		input  exception_t                      lsu_exception_o,  // address translation threw an exception //output
		// General control signals
		input riscv::priv_lvl_t                 priv_lvl_i,
		input riscv::priv_lvl_t                 ld_st_priv_lvl_i,
		input logic                             sum_i,
		input logic                             mxr_i,
		// input logic flag_mprv_i,
		input logic [riscv::PPNW-1:0]           satp_ppn_i,
		input logic [ASID_WIDTH-1:0]            asid_i,
		input logic [ASID_WIDTH-1:0]            asid_to_be_flushed_i,
		input logic [riscv::VLEN-1:0]           vaddr_to_be_flushed_i,
		input logic                             flush_tlb_i,
		// Performance counters
		input  logic                            itlb_miss_o, //output
		input  logic                            dtlb_miss_o, //output
		// PTW memory interface
		input  dcache_req_o_t                   req_port_i,
		input  dcache_req_i_t                   req_port_o, //output
		// PMP
		input  riscv::pmpcfg_t [15:0]           pmpcfg_i,
		input  logic [15:0][riscv::PLEN-1:0]    pmpaddr_i
	);

//==============================================================================
// Local Parameters
//==============================================================================

genvar j;
default clocking cb @(posedge clk_i);
endclocking
default disable iff (!rst_ni);
reg reset_r = 0;
am__rst: assume property (reset_r != !rst_ni);
always_ff @(posedge clk_i)
    reset_r <= 1'b1;

// Re-defined wires 
wire itlb_req_val;
wire itlb_req_rdy;
wire [riscv::VLEN+ASID_WIDTH-1:0] itlb_req_stable;
wire itlb_res_val;
wire dtlb_req_val;
wire [riscv::VLEN+ASID_WIDTH-1:0] dtlb_req_stable;
wire dtlb_res_val;

// Symbolics and Handshake signals
wire dtlb_res_hsk = dtlb_res_val;
wire dtlb_req_hsk = dtlb_req_val;
wire itlb_res_hsk = itlb_res_val;
wire itlb_req_hsk = itlb_req_val && itlb_req_rdy;

//==============================================================================
// Modeling
//==============================================================================

// Modeling incoming request for dtlb_lookup
// Generate sampling signals and model
reg [3:0] dtlb_lookup_transid_sampled;
wire dtlb_lookup_transid_set = dtlb_req_hsk;
wire dtlb_lookup_transid_response = dtlb_res_hsk;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		dtlb_lookup_transid_sampled <= '0;
	end else if (dtlb_lookup_transid_set || dtlb_lookup_transid_response ) begin
		dtlb_lookup_transid_sampled <= dtlb_lookup_transid_sampled + dtlb_lookup_transid_set - dtlb_lookup_transid_response;
	end
end
co__dtlb_lookup_transid_sampled: cover property (|dtlb_lookup_transid_sampled);
if (ASSERT_INPUTS) begin
	as__dtlb_lookup_transid_sample_no_overflow: assert property (dtlb_lookup_transid_sampled != '1 || !dtlb_lookup_transid_set);
end else begin
	am__dtlb_lookup_transid_sample_no_overflow: assume property (dtlb_lookup_transid_sampled != '1 || !dtlb_lookup_transid_set);
end


// Assert that every request has a response and that every reponse has a request
as__dtlb_lookup_transid_eventual_response: assert property (dtlb_lookup_transid_set |-> s_eventually(dtlb_res_val));
as__dtlb_lookup_transid_was_a_request: assert property (dtlb_lookup_transid_response |-> dtlb_lookup_transid_set || dtlb_lookup_transid_sampled);

// Modeling incoming request for itlb_lookup
// Generate sampling signals and model
reg [3:0] itlb_lookup_transid_sampled;
wire itlb_lookup_transid_set = itlb_req_hsk;
wire itlb_lookup_transid_response = itlb_res_hsk;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		itlb_lookup_transid_sampled <= '0;
	end else if (itlb_lookup_transid_set || itlb_lookup_transid_response ) begin
		itlb_lookup_transid_sampled <= itlb_lookup_transid_sampled + itlb_lookup_transid_set - itlb_lookup_transid_response;
	end
end
if (ASSERT_INPUTS) begin
	as__itlb_lookup_transid_sample_no_overflow: assert property (itlb_lookup_transid_sampled != '1 || !itlb_lookup_transid_set);
end else begin
	am__itlb_lookup_transid_sample_no_overflow: assume property (itlb_lookup_transid_sampled != '1 || !itlb_lookup_transid_set);
end


// Assume payload is stable and valid is non-dropping
if (ASSERT_INPUTS) begin
	as__itlb_lookup_transid_stability: assert property (itlb_req_val && !itlb_req_rdy |=> itlb_req_val && $stable(itlb_req_stable) );
end else begin
	am__itlb_lookup_transid_stability: assume property (itlb_req_val && !itlb_req_rdy |=> itlb_req_val && $stable(itlb_req_stable) );
end

// Assert that if valid eventually ready or dropped valid
as__itlb_lookup_transid_hsk_or_drop: assert property (itlb_req_val |-> s_eventually(!itlb_req_val || itlb_req_rdy));
// Assert that every request has a response and that every reponse has a request
as__itlb_lookup_transid_eventual_response: assert property (itlb_lookup_transid_set |-> s_eventually(itlb_res_val));
as__itlb_lookup_transid_was_a_request: assert property (itlb_lookup_transid_response |-> itlb_lookup_transid_set || itlb_lookup_transid_sampled);

assign itlb_res_val = icache_areq_o.fetch_valid;
assign itlb_req_stable = {asid_i,icache_areq_i.fetch_vaddr};
assign itlb_req_rdy = icache_areq_o.fetch_valid;
assign dtlb_req_stable = {asid_i, lsu_vaddr_i};
assign itlb_req_val = icache_areq_i.fetch_req;
assign dtlb_res_val = lsu_valid_o;
assign dtlb_req_val = lsu_req_i;

//X PROPAGATION ASSERTIONS
`ifdef XPROP
	 as__no_x_itlb_req_val: assert property(!$isunknown(itlb_req_val));
	 as__no_x_itlb_req_stable: assert property(itlb_req_val |-> !$isunknown(itlb_req_stable));
	 as__no_x_dtlb_req_val: assert property(!$isunknown(dtlb_req_val));
	 as__no_x_dtlb_req_stable: assert property(dtlb_req_val |-> !$isunknown(dtlb_req_stable));
`endif

//====DESIGNER-ADDED-SVA====//
//Assume inputs (vaddr and asid) are stable while transaction not satisfied
am__itrans : assume property (enable_translation_i);
am__dtrans : assume property (en_ld_st_translation_i);
am__no_flush : assume property (!flush_i);
am__no_flush_itlb : assume property (!flush_tlb_i);
am__no_dtlb_forever: assume property (dtlb_req_hsk |=> s_eventually(!dtlb_req_val));
endmodule