// The Clear BSD License
// Copyright (c) [2021] [The Trustees of Princeton University]
// All rights reserved.
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted for academic and research use only (subject to the 
// limitations in the disclaimer below) provided that the following conditions are met:
//     * Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
// 
//     * Redistributions in binary form must reproduce the above copyright
//     notice, this list of conditions and the following disclaimer in the
//     documentation and/or other materials provided with the distribution.
// 
//     * Neither the name of the copyright holder nor the names of its
//     contributors may be used to endorse or promote products derived from this
//     software without specific prior written permission.
// 
// NO EXPRESS OR IMPLIED LICENSES TO ANY PARTY'S PATENT RIGHTS ARE GRANTED BY
// THIS LICENSE. THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND
// CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
// PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
// CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,
// EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
// PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
// IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
// 
// This property file was autogenerated by AutoSVA on 2021-04-06
// to check the behavior of the original RTL module, whose interface is described below: 


module tlb_prop
 import ariane_pkg::*; #(
		parameter ASSERT_INPUTS = 0,
		parameter int unsigned TLB_ENTRIES = 4,
		parameter int unsigned ASID_WIDTH  = 1
)(
		input  logic                    clk_i,    // Clock
		input  logic                    rst_ni,   // Asynchronous reset active low
		input  logic                    flush_i,  // Flush signal
		// Update TLB
		input  tlb_update_t             update_i,
		// Lookup signals
		input  logic                    lu_access_i,
		input  logic [ASID_WIDTH-1:0]   lu_asid_i,
		input  logic [riscv::VLEN-1:0]  lu_vaddr_i,
		input  riscv::pte_t             lu_content_o, //output
		input  logic [ASID_WIDTH-1:0]   asid_to_be_flushed_i,
		input  logic [riscv::VLEN-1:0]  vaddr_to_be_flushed_i,
		input  logic                    lu_is_2M_o, //output
		input  logic                    lu_is_1G_o, //output
		input  logic                    lu_hit_o //output
	);

//==============================================================================
// Local Parameters
//==============================================================================

genvar j;
default clocking cb @(posedge clk_i);
endclocking
default disable iff (!rst_ni);
reg reset_r = 0;
am__rst: assume property (reset_r != !rst_ni);
always_ff @(posedge clk_i)
    reset_r <= 1'b1;

// Re-defined wires 
wire lk_req_val;
wire lk_req_rdy;
wire [riscv::VLEN+ASID_WIDTH-1:0] lk_req_stable;
wire lk_res_val;
wire miss_val;
wire [27:0] miss_data;
wire alloc_val;
wire [27:0] alloc_data;

// Symbolics and Handshake signals
wire lk_res_hsk = lk_res_val;
wire lk_req_hsk = lk_req_val && lk_req_rdy;
wire alloc_hsk = alloc_val;
wire miss_hsk = miss_val;

//==============================================================================
// Modeling
//==============================================================================

// Modeling incoming request for lookup
// Generate sampling signals and model
reg [3:0] lookup_transid_sampled;
wire lookup_transid_set = lk_req_hsk;
wire lookup_transid_response = lk_res_hsk;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		lookup_transid_sampled <= '0;
	end else if (lookup_transid_set || lookup_transid_response ) begin
		lookup_transid_sampled <= lookup_transid_sampled + lookup_transid_set - lookup_transid_response;
	end
end
if (ASSERT_INPUTS) begin
	as__lookup_transid_sample_no_overflow: assert property (lookup_transid_sampled != '1 || !lookup_transid_set);
end else begin
	am__lookup_transid_sample_no_overflow: assume property (lookup_transid_sampled != '1 || !lookup_transid_set);
end


// Assume payload is stable and valid is non-dropping
if (ASSERT_INPUTS) begin
	as__lookup_transid_stability: assert property (lk_req_val && !lk_req_rdy |=> lk_req_val && $stable(lk_req_stable) );
end else begin
	am__lookup_transid_stability: assume property (lk_req_val && !lk_req_rdy |=> lk_req_val && $stable(lk_req_stable) );
end

// Assert that if valid eventually ready or dropped valid
as__lookup_transid_hsk_or_drop: assert property (lk_req_val |-> s_eventually(!lk_req_val || lk_req_rdy));
// Assert that every request has a response and that every reponse has a request
as__lookup_transid_eventual_response: assert property (lookup_transid_set |-> s_eventually(lk_res_val));
as__lookup_transid_was_a_request: assert property (lookup_transid_response |-> lookup_transid_set || lookup_transid_sampled);

// Modeling outstanding request for update
reg [1-1:0] update_outstanding_req_r;
reg [1-1:0][27:0] update_outstanding_req_data_r;

always_ff @(posedge clk_i) begin
	if(!rst_ni) begin
		update_outstanding_req_r <= '0;
	end else begin
		if (miss_hsk) begin
			update_outstanding_req_r <= 1'b1;
			update_outstanding_req_data_r <= miss_data;
		end
		if (alloc_hsk) begin
			update_outstanding_req_r <= 1'b0;
		end
	end
end


generate
if (ASSERT_INPUTS) begin : update_gen
	as__update1: assert property (!update_outstanding_req_r |-> !(alloc_hsk));
	as__update2: assert property (update_outstanding_req_r |-> s_eventually(alloc_hsk&&
	 (alloc_data == update_outstanding_req_data_r) ));
end else begin : update_else_gen
	for ( j = 0; j < 1; j = j + 1) begin : update_for_gen
		co__update: cover property (update_outstanding_req_r[j]);
		am__update1: assume property (!update_outstanding_req_r[j] |-> !(alloc_val));
		am__update2: assume property (update_outstanding_req_r[j] |-> s_eventually(alloc_val&&
	 (alloc_data == update_outstanding_req_data_r[j]) ));
	end
end
endgenerate

assign alloc_data = {update_i.asid,update_i.vpn};
assign lk_req_stable = {lu_vaddr_i, lu_asid_i};
assign miss_val = lu_access_i && !lu_hit_o;
assign alloc_val = update_i.valid;
assign lk_res_val = lu_access_i && lu_hit_o;
assign lk_req_rdy = lu_access_i && lu_hit_o;
assign lk_req_val = lu_access_i;
assign miss_data = {lu_asid_i,lu_vaddr_i[38:12]};

//X PROPAGATION ASSERTIONS
`ifdef XPROP
	 as__no_x_miss_val: assert property(!$isunknown(miss_val));
	 as__no_x_miss_data: assert property(miss_val |-> !$isunknown(miss_data));
	 as__no_x_alloc_val: assert property(!$isunknown(alloc_val));
	 as__no_x_alloc_data: assert property(alloc_val |-> !$isunknown(alloc_data));
	 as__no_x_lk_req_val: assert property(!$isunknown(lk_req_val));
	 as__no_x_lk_req_stable: assert property(lk_req_val |-> !$isunknown(lk_req_stable));
`endif

//====DESIGNER-ADDED-SVA====//
am__no_flush: assume property (flush_i=='0);
endmodule