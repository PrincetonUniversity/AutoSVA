bind tlb tlb_prop
	#(
		.ASSERT_INPUTS (0)
	) u_tlb_sva(.*);